// ======================================================================
// Affiliation:			Tsinghua Univ
// Author:				Yongxiang Guo
// Create Date:			Oct 23, 2022
// Module Name:			decoder1
// Description:			full subtractor
// Additional Comments:	VL17 on nowcoder
// ======================================================================

`timescale 1ns/1ns

module decoder1 (
	input	wire				A,
	input	wire				B,
	input	wire				Ci,
	output	wire				D,
	output	wire				Co
);

wire	Y0n;
wire	Y1n;
wire	Y2n;
wire	Y3n;
wire	Y4n;
wire	Y5n;
wire	Y6n;
wire	Y7n;

//			A	B	Ci		D	Co
//	Y0n		0	0	0		0	0
//	Y1n		0	0	1		1	1
//	Y2n		0	1	0		1	1
//	Y3n		0	1	1		0	1
//	Y4n		1	0	0		1	0
//	Y5n		1	0	1		0	0
//	Y6n		1	1	0		0	0
//	Y7n		1	1	1		1	1
assign D  = ~(Y1n & Y2n & Y4n & Y7n);
assign Co = ~(Y1n & Y2n & Y3n & Y7n);

decoder_38 u_decoder_38(
	.E 			( 1'b1 ),
	.A0			( Ci   ),
	.A1			( B    ),
	.A2			( A    ),

	.Y0n		( Y0n  ),  
	.Y1n		( Y1n  ), 
	.Y2n		( Y2n  ), 
	.Y3n		( Y3n  ), 
	.Y4n		( Y4n  ), 
	.Y5n		( Y5n  ), 
	.Y6n		( Y6n  ), 
	.Y7n		( Y7n  )
);

endmodule


module decoder_38(
   input             E      ,
   input             A0     ,
   input             A1     ,
   input             A2     ,
   
   output reg       Y0n    ,  
   output reg       Y1n    , 
   output reg       Y2n    , 
   output reg       Y3n    , 
   output reg       Y4n    , 
   output reg       Y5n    , 
   output reg       Y6n    , 
   output reg       Y7n    
);

always @(*)begin
   if(!E)begin
      Y0n = 1'b1;
      Y1n = 1'b1;
      Y2n = 1'b1;
      Y3n = 1'b1;
      Y4n = 1'b1;
      Y5n = 1'b1;
      Y6n = 1'b1;
      Y7n = 1'b1;
   end  
   else begin
      case({A2,A1,A0})
         3'b000 : begin
                     Y0n = 1'b0; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b1;
                  end 
         3'b001 : begin
                     Y0n = 1'b1; Y1n = 1'b0; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b1;
                  end 
         3'b010 : begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b0; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b1;
                  end 
         3'b011 : begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b0; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b1;
                  end 
         3'b100 : begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b0; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b1;
                  end 
         3'b101 : begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b0; Y6n = 1'b1; Y7n = 1'b1;
                  end 
         3'b110 : begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b0; Y7n = 1'b1;
                  end 
         3'b111 : begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b0;
                  end 
         default: begin
                     Y0n = 1'b1; Y1n = 1'b1; Y2n = 1'b1; Y3n = 1'b1; 
                     Y4n = 1'b1; Y5n = 1'b1; Y6n = 1'b1; Y7n = 1'b1;
                  end
      endcase  
   end 
end    
     
endmodule

