// ======================================================================
// Copyright (c) 2023-2023 All rights reserved
// ======================================================================
// Affiliation  : Tsinghua Univ & NeuraMatrix
// Author       : Yongxiang Guo
// Create Date  : 2023-06-09 13:34:00
// Revise Date  : 2023-06-09 13:34:02
// File Name    : sfifo.v
// Description  : VL68 on nowcoder
// ======================================================================

module dual_port_RAM #(
  parameter DEPTH = 16,
  parameter WIDTH = 8
) (
  input  wire                     wclk,
  input  wire                     wenc,
  input  wire [$clog2(DEPTH)-1:0] waddr,
  input  wire [WIDTH-1:0]         wdata,
  input  wire                     rclk,
  input  wire                     renc,
  input  wire [$clog2(DEPTH)-1:0] raddr,
  output reg  [WIDTH-1:0]         rdata
);

  reg [WIDTH-1:0] RAM_MEM [0:DEPTH-1];

  always @(posedge wclk) begin
    if(wenc)
      RAM_MEM[waddr] <= wdata;
  end

  always @(posedge rclk) begin
    if(renc)
      rdata <= RAM_MEM[raddr];
  end

endmodule


module sfifo #(
  parameter WIDTH = 8,
  parameter DEPTH = 16
)(
  input  wire             clk   ,
  input  wire             rst_n ,
  input  wire             winc  ,
  input  wire             rinc  ,
  input  wire [WIDTH-1:0] wdata ,

  output wire             wfull ,
  output wire             rempty,
  output wire [WIDTH-1:0] rdata
);

  localparam ADDR_WIDTH = $clog2(DEPTH);

  wire [ADDR_WIDTH-1:0] waddr;
  wire [ADDR_WIDTH-1:0] raddr;
  wire                  renc;
  wire                  wenc;
  wire                  full;
  wire                  empty;

  reg  [ADDR_WIDTH:0]   waddr_reg;
  reg  [ADDR_WIDTH:0]   raddr_reg;
  reg                   full_reg;
  reg                   empty_reg;

  assign waddr = waddr_reg[ADDR_WIDTH-1:0];
  assign raddr = raddr_reg[ADDR_WIDTH-1:0];
  assign wenc = winc & (~full);
  assign renc = rinc & (~empty);

  // Write fifo
  always @(posedge clk or negedge rst_n) begin
    if (~rst_n) begin
      waddr_reg <= {(ADDR_WIDTH+1){1'b0}};
    end else begin
      if (wenc) begin
        if (waddr_reg == DEPTH - 1) begin
          waddr_reg[ADDR_WIDTH-1:0] <= {ADDR_WIDTH{1'b0}};
          waddr_reg[ADDR_WIDTH] <= ~waddr_reg[ADDR_WIDTH];
        end else begin
          waddr_reg <= waddr_reg + 1'd1;
        end
      end
    end
  end

  // Read fifo
  always @(posedge clk or negedge rst_n) begin
    if (~rst_n) begin
      raddr_reg <= {(ADDR_WIDTH+1){1'b0}};
    end else begin
      if (renc) begin
        if (raddr_reg == DEPTH - 1) begin
          raddr_reg[ADDR_WIDTH-1:0] <= {ADDR_WIDTH{1'b0}};
          raddr_reg[ADDR_WIDTH] <= ~raddr_reg[ADDR_WIDTH];
        end else begin
          raddr_reg <= raddr_reg + 1'd1;
        end
      end
    end
  end

  // Full flag
  // Nowcoder answer is wrong
  assign full = ({~waddr_reg[ADDR_WIDTH], waddr_reg[ADDR_WIDTH-1:0]} == raddr_reg) ? 1'b1 : 1'b0;
  always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
      full_reg <= 1'b0;
    end else begin
      full_reg <= full;
    end
  end
  assign wfull = full_reg;
  // This is the right logic: wfull should not delay 1 cycle
  // assign wfull = ({~waddr_reg[ADDR_WIDTH], waddr_reg[ADDR_WIDTH-1:0]} == raddr_reg) ? 1'b1 : 1'b0;

  // Empty flag
  // Nowcoder answer is wrong
  assign empty = (waddr_reg == raddr_reg) ? 1'b1 : 1'b0;
  always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
      empty_reg <= 1'b0;
    end else begin
      empty_reg <= empty;
    end
  end
  assign rempty = empty_reg;
  // This is the right logic: rempty should not delay 1 cycle
  // assign rempty = (waddr_reg == raddr_reg) ? 1'b1 : 1'b0;

  dual_port_RAM #(
    .DEPTH ( DEPTH ),
    .WIDTH ( WIDTH )
  ) i_dual_port_RAM (
    .wclk  ( clk   ),
    .wenc  ( wenc  ),
    .waddr ( waddr ),
    .wdata ( wdata ),
    .rclk  ( clk   ),
    .renc  ( renc  ),
    .raddr ( raddr ),
    .rdata ( rdata )
  );

endmodule